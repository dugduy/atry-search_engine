{"name": "c.SV"}