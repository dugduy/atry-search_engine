{"name": "d.SV"}