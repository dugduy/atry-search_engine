{"name": "b.SV", "title": "Site Yap\u0131m A\u015famas\u0131ndad\u0131r"}